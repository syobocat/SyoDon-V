module httpsig

//import crypto.ed25519
//import crypto.pem
//import crypto.sha512
//import encoding.base64
//import net.http
//import user

pub fn verify_header() ! {
	// TODO
}
