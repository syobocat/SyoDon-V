module httpsig

//import crypto.ed25519
//import crypto.pem
//import crypto.sha256
//import crypto.sha512
//import encoding.base64
//import user

pub fn verify_headers_rfc9421(params HttpsigInput) ! {
	// TODO
}
